 
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2distance IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;    
--		Switch			: 	in		std_logic;		
      v_in        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      distance       :  OUT   STD_LOGIC_VECTOR(12 DOWNTO 0));

END voltage2distance;

ARCHITECTURE behavior OF voltage2distance IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.
-- See how to get the distance output at the bottom of this file,
-- after begin.

type array_1d is array (0 to 4095) of integer;
constant v2d_far : array_1d := (

(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	3296	)	,
(	3288	)	,
(	3279	)	,
(	3270	)	,
(	3262	)	,
(	3253	)	,
(	3245	)	,
(	3237	)	,
(	3228	)	,
(	3220	)	,
(	3212	)	,
(	3203	)	,
(	3195	)	,
(	3187	)	,
(	3179	)	,
(	3171	)	,
(	3163	)	,
(	3155	)	,
(	3147	)	,
(	3139	)	,
(	3131	)	,
(	3123	)	,
(	3116	)	,
(	3108	)	,
(	3100	)	,
(	3093	)	,
(	3085	)	,
(	3077	)	,
(	3070	)	,
(	3062	)	,
(	3055	)	,
(	3047	)	,
(	3040	)	,
(	3032	)	,
(	3025	)	,
(	3018	)	,
(	3011	)	,
(	3003	)	,
(	2996	)	,
(	2989	)	,
(	2982	)	,
(	2975	)	,
(	2968	)	,
(	2961	)	,
(	2953	)	,
(	2947	)	,
(	2940	)	,
(	2933	)	,
(	2926	)	,
(	2919	)	,
(	2912	)	,
(	2905	)	,
(	2899	)	,
(	2892	)	,
(	2885	)	,
(	2878	)	,
(	2872	)	,
(	2865	)	,
(	2859	)	,
(	2852	)	,
(	2846	)	,
(	2839	)	,
(	2833	)	,
(	2826	)	,
(	2820	)	,
(	2813	)	,
(	2807	)	,
(	2801	)	,
(	2794	)	,
(	2788	)	,
(	2782	)	,
(	2776	)	,
(	2770	)	,
(	2763	)	,
(	2757	)	,
(	2751	)	,
(	2745	)	,
(	2739	)	,
(	2733	)	,
(	2727	)	,
(	2721	)	,
(	2715	)	,
(	2709	)	,
(	2703	)	,
(	2697	)	,
(	2692	)	,
(	2686	)	,
(	2680	)	,
(	2674	)	,
(	2668	)	,
(	2663	)	,
(	2657	)	,
(	2651	)	,
(	2646	)	,
(	2640	)	,
(	2634	)	,
(	2629	)	,
(	2623	)	,
(	2618	)	,
(	2612	)	,
(	2607	)	,
(	2601	)	,
(	2596	)	,
(	2590	)	,
(	2585	)	,
(	2580	)	,
(	2574	)	,
(	2569	)	,
(	2564	)	,
(	2558	)	,
(	2553	)	,
(	2548	)	,
(	2543	)	,
(	2537	)	,
(	2532	)	,
(	2527	)	,
(	2522	)	,
(	2517	)	,
(	2512	)	,
(	2507	)	,
(	2501	)	,
(	2496	)	,
(	2491	)	,
(	2486	)	,
(	2481	)	,
(	2476	)	,
(	2471	)	,
(	2467	)	,
(	2462	)	,
(	2457	)	,
(	2452	)	,
(	2447	)	,
(	2442	)	,
(	2437	)	,
(	2433	)	,
(	2428	)	,
(	2423	)	,
(	2418	)	,
(	2414	)	,
(	2409	)	,
(	2404	)	,
(	2399	)	,
(	2395	)	,
(	2390	)	,
(	2386	)	,
(	2381	)	,
(	2376	)	,
(	2372	)	,
(	2367	)	,
(	2363	)	,
(	2358	)	,
(	2354	)	,
(	2349	)	,
(	2345	)	,
(	2340	)	,
(	2336	)	,
(	2332	)	,
(	2327	)	,
(	2323	)	,
(	2318	)	,
(	2314	)	,
(	2310	)	,
(	2305	)	,
(	2301	)	,
(	2297	)	,
(	2293	)	,
(	2288	)	,
(	2284	)	,
(	2280	)	,
(	2276	)	,
(	2271	)	,
(	2267	)	,
(	2263	)	,
(	2259	)	,
(	2255	)	,
(	2251	)	,
(	2247	)	,
(	2242	)	,
(	2238	)	,
(	2234	)	,
(	2230	)	,
(	2226	)	,
(	2222	)	,
(	2218	)	,
(	2214	)	,
(	2210	)	,
(	2206	)	,
(	2202	)	,
(	2198	)	,
(	2194	)	,
(	2191	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2175	)	,
(	2171	)	,
(	2167	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2148	)	,
(	2145	)	,
(	2141	)	,
(	2137	)	,
(	2134	)	,
(	2130	)	,
(	2126	)	,
(	2122	)	,
(	2119	)	,
(	2115	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2101	)	,
(	2097	)	,
(	2094	)	,
(	2090	)	,
(	2086	)	,
(	2083	)	,
(	2079	)	,
(	2076	)	,
(	2072	)	,
(	2069	)	,
(	2065	)	,
(	2062	)	,
(	2058	)	,
(	2055	)	,
(	2052	)	,
(	2048	)	,
(	2045	)	,
(	2041	)	,
(	2038	)	,
(	2035	)	,
(	2031	)	,
(	2028	)	,
(	2024	)	,
(	2021	)	,
(	2018	)	,
(	2014	)	,
(	2011	)	,
(	2008	)	,
(	2005	)	,
(	2001	)	,
(	1998	)	,
(	1995	)	,
(	1992	)	,
(	1988	)	,
(	1985	)	,
(	1982	)	,
(	1979	)	,
(	1975	)	,
(	1972	)	,
(	1969	)	,
(	1966	)	,
(	1963	)	,
(	1960	)	,
(	1957	)	,
(	1953	)	,
(	1950	)	,
(	1947	)	,
(	1944	)	,
(	1941	)	,
(	1938	)	,
(	1935	)	,
(	1932	)	,
(	1929	)	,
(	1926	)	,
(	1923	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1908	)	,
(	1905	)	,
(	1902	)	,
(	1899	)	,
(	1896	)	,
(	1893	)	,
(	1890	)	,
(	1887	)	,
(	1884	)	,
(	1881	)	,
(	1878	)	,
(	1876	)	,
(	1873	)	,
(	1870	)	,
(	1867	)	,
(	1864	)	,
(	1861	)	,
(	1858	)	,
(	1856	)	,
(	1853	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1842	)	,
(	1839	)	,
(	1836	)	,
(	1833	)	,
(	1831	)	,
(	1828	)	,
(	1825	)	,
(	1822	)	,
(	1820	)	,
(	1817	)	,
(	1814	)	,
(	1812	)	,
(	1809	)	,
(	1806	)	,
(	1803	)	,
(	1801	)	,
(	1798	)	,
(	1796	)	,
(	1793	)	,
(	1790	)	,
(	1788	)	,
(	1785	)	,
(	1782	)	,
(	1780	)	,
(	1777	)	,
(	1775	)	,
(	1772	)	,
(	1769	)	,
(	1767	)	,
(	1764	)	,
(	1762	)	,
(	1759	)	,
(	1757	)	,
(	1754	)	,
(	1752	)	,
(	1749	)	,
(	1747	)	,
(	1744	)	,
(	1742	)	,
(	1739	)	,
(	1737	)	,
(	1734	)	,
(	1732	)	,
(	1729	)	,
(	1727	)	,
(	1724	)	,
(	1722	)	,
(	1719	)	,
(	1717	)	,
(	1715	)	,
(	1712	)	,
(	1710	)	,
(	1707	)	,
(	1705	)	,
(	1703	)	,
(	1700	)	,
(	1698	)	,
(	1696	)	,
(	1693	)	,
(	1691	)	,
(	1688	)	,
(	1686	)	,
(	1684	)	,
(	1681	)	,
(	1679	)	,
(	1677	)	,
(	1674	)	,
(	1672	)	,
(	1670	)	,
(	1668	)	,
(	1665	)	,
(	1663	)	,
(	1661	)	,
(	1658	)	,
(	1656	)	,
(	1654	)	,
(	1652	)	,
(	1649	)	,
(	1647	)	,
(	1645	)	,
(	1643	)	,
(	1641	)	,
(	1638	)	,
(	1636	)	,
(	1634	)	,
(	1632	)	,
(	1630	)	,
(	1627	)	,
(	1625	)	,
(	1623	)	,
(	1621	)	,
(	1619	)	,
(	1617	)	,
(	1614	)	,
(	1612	)	,
(	1610	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1602	)	,
(	1599	)	,
(	1597	)	,
(	1595	)	,
(	1593	)	,
(	1591	)	,
(	1589	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1581	)	,
(	1579	)	,
(	1577	)	,
(	1575	)	,
(	1573	)	,
(	1570	)	,
(	1568	)	,
(	1566	)	,
(	1564	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1552	)	,
(	1550	)	,
(	1548	)	,
(	1546	)	,
(	1544	)	,
(	1542	)	,
(	1541	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1533	)	,
(	1531	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1517	)	,
(	1515	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1499	)	,
(	1497	)	,
(	1495	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1480	)	,
(	1478	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1468	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1447	)	,
(	1445	)	,
(	1443	)	,
(	1441	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1423	)	,
(	1421	)	,
(	1419	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1403	)	,
(	1401	)	,
(	1400	)	,
(	1398	)	,
(	1396	)	,
(	1395	)	,
(	1393	)	,
(	1391	)	,
(	1390	)	,
(	1388	)	,
(	1387	)	,
(	1385	)	,
(	1383	)	,
(	1382	)	,
(	1380	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1374	)	,
(	1372	)	,
(	1371	)	,
(	1369	)	,
(	1368	)	,
(	1366	)	,
(	1365	)	,
(	1363	)	,
(	1362	)	,
(	1360	)	,
(	1359	)	,
(	1357	)	,
(	1355	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1349	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1339	)	,
(	1337	)	,
(	1336	)	,
(	1334	)	,
(	1333	)	,
(	1331	)	,
(	1330	)	,
(	1329	)	,
(	1327	)	,
(	1326	)	,
(	1324	)	,
(	1323	)	,
(	1321	)	,
(	1320	)	,
(	1318	)	,
(	1317	)	,
(	1315	)	,
(	1314	)	,
(	1313	)	,
(	1311	)	,
(	1310	)	,
(	1308	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1303	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1285	)	,
(	1283	)	,
(	1282	)	,
(	1280	)	,
(	1279	)	,
(	1278	)	,
(	1276	)	,
(	1275	)	,
(	1274	)	,
(	1272	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1266	)	,
(	1264	)	,
(	1263	)	,
(	1262	)	,
(	1260	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1241	)	,
(	1239	)	,
(	1238	)	,
(	1237	)	,
(	1236	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1231	)	,
(	1229	)	,
(	1228	)	,
(	1227	)	,
(	1225	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1220	)	,
(	1219	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1209	)	,
(	1208	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	287	)	
);



--constant v2d_close : array_1d := (
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	100	)	,
--(	200	)	,
--(	300	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	,
--(	0	)	
--);

begin
   -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
	distance <= std_logic_vector(to_unsigned(v2d_far(to_integer(unsigned(v_in))),distance'length));
--				process (switch, clk)
--					begin	
--					if	rising_edge(clk) then
--						if			Switch ='0' then
--							distance <= std_logic_vector(to_unsigned(v2d_far(to_integer(unsigned(voltage))),distance'length));
--						elsif 	Switch ='1' then
--							distance <= std_logic_vector(to_unsigned(v2d_close(to_integer(unsigned(voltage))),distance'length));
--						end if;
--					end if;	
--				end process; 	
--   

end behavior;
